19D070052 Sheel Shah Expt3 CE Amp Biasing
.model bc547a NPN IS=10f BF=400 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f
** nodes:
**   1 Vin, 2 Rs-C1, 3 base1
**   4 emitter1
**   5 collector1, 6 base2
**   7 emitter2, 8 Re2    
**   9 vcc/collector2
**   10 vout
vin 1 0 dc 0 ac 10m
vcc 9 0 12

rs 1 2 0
c1 2 3 10u

q1 5 3 4 bc547a
r2 3 0 2.2k
r1 3 9 10k
re 4 0 1k
ce 4 0 100u
rc 5 9 1.2k

vib2 5 6 0
vie2 7 8 0

q2 9 6 7 bc547a
re2 8 0 10k
c2 7 10 10u
rl 10 0 10k

.op
.control
run
print i(vib2) i(vie2)
.endc
.end
