Sheel Shah 19D070052 Expt4 Diff Pair

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

** nodes:
** 1 emitter of both
** 2 base1, 3 base2
** 20 in1, 30 in2
** 4 collector1, 5 collector2
** 6 vee, 7 vcc
q1 4 2 1 bc547a
q2 5 3 1 bc547a

v_cc 7 0 12
v_ic1 7 74 0
r_c1 74 4 6.8k
v_ic2 7 75 0
r_c2 75 5 6.8k

v_i1 20 0
r_b1 2 20 1k
v_i2 30 0 0
r_b2 3 30 1k

v_ee 6 0 -12
r_e 6 1 10k

.dc v_i1 -1 1 0.1
.control
run
plot v(4), v(5)
.endc
.end