Sheel Shah 19D070052 Expt4 Current Source

.include all_model_files/zener_B.txt
.model bc557a PNP IS=10f BF=100 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

** nodes:
** 1 vcc, 2 emitter, 3 base, 4/5 collector
q1 4 3 2 bc557a
v_cc 1 0 12
x_z 3 1 DI_1N4734A
r_e 1 2 4.7k
r_b 3 0 2.2k
v0 4 5 0
r_l 5 0 1k

.op
.control
run
print v(2), v(3), v(4), i(v0)
.endc
.end
