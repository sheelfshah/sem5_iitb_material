Sheel Shah 19D070052 Expt4 Current Mirror

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f

** nodes:
** 1 vcc
** 2 collector1/base1/base2
** 3 collector2/vout
q1 2 2 0 bc547a
q2 3 2 0 bc547a
v_cc 1 0 12
v_out 3 0 1
r0 1 2 10k

.op
.control
run
print i(v_out), i(v_cc), v(2)
.endc
.end