Integrator
.include all_model_files/ua741.txt

* describe circuit
* <element name> <nodes list> <value>
* voltage_nodename positive_node negative_node dc_value/function
    * v 1 0 5
* sine voltage: sin(offset amplitude frequency time_delay damping_factor)
    * v 1 0 sin(0 2 1k 0 0)
* peicewise linear: pwl(time1 value1 time2 value2 ...)
    * v 1 0 pwl(0 0 10m 0 11m 5 20m 5)
* pulse waveform: pulse(initial-value pulsed-value TD TR TF PW period)
    * v 1 0 pulse(0 1 1m 1m 1m 6m 10m)
* exponentioal waveform: exp(initial pulsed rise-delay rise-time fall-delay fall-time)
    * v 1 0 exp(1 0 10m 10m 10m 10m)
* ac analysis: dc dc_val ac ac_val
    * v 1 0 dc 0 ac 1
x0 0 1 2 3 4 ua741
r0 5 1 1k
c0 4 1 0.1u
v1 2 0 15
v2 3 0 -15
v0 5 0 sin(0 2 1k 0 0)


* dc analysis: dc node_name initial_value final_value step
    * .dc v 0 5 0.1
* transient analysis: tran timestep end_time
    * .tran 10u 20m
* ac analysis: ac lin/dec num_points start_freq end_freq
    * .ac dec 10 1 1k
.tran 20u 12m

* start control
.control

run

* plot vdb(2); plots magnitude in dB
* plot phase(v(2)); plots phase of v(2)
* plot i(v); plots current through voltage_element v, only voltage elements allowed
* plot v(1) vs v(2); for output vs input
* use dummy voltage elements to measure current through all elements
plot v(5) vs v(4)

* hardcopy filename.ps plotting_value

* end control
.endc

.end